systemverilog information is here
