systemverilog information is not here
write something into sys.sv
do something change
<<<<<<< HEAD
create  a new branch is quick & simple
=======
add a newbranch is quick and simple.

>>>>>>> feature1

ajjdhhd
abvcckkcl
