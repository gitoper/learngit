jkfskjfksjsk
