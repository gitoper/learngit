systemverilog information is here
write something into sys.sv
do something change
add a newbranch is quick AND simple.

