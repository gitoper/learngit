systemverilog information is here
write something into sys.sv
do something change
create  a new branch is quick & simple
