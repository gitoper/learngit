adkdhakdhal
