systemverilog information is here
write something into sys.sv
do something change
