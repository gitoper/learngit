systemverilog information is here
write something into sys.sv
